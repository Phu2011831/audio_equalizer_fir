library verilog;
use verilog.vl_types.all;
entity audio_equalizer_tb is
end audio_equalizer_tb;
