//module audio_equalizer_tb();
