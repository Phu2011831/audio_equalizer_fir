`timescale 1ns / 1ps

`ifndef CONSTANTS
`define CONSTANTS

	`define ORDER_FIR 		64
	`define GAIN_BAND_1		5'd9
	`define GIAN_BAND_2		5'd8
	`define GIAN_BAND_3		5'd7
	`define GIAN_BAND_4		5'd6
	`define GIAN_BAND_5		5'd5
	`define GIAN_BAND_6		5'd4
	`define GIAN_BAND_7		5'd3
	`define GIAN_BAND_8		5'd2
	`define GIAN_BAND_9		5'd1
	`define INPUT_WIDTH		24
	`define OUTPUT_WIDTH		24
	`define NUMBER_BANDS		9



`endif